// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 15.0.0 Build 145 04/22/2015 SJ Web Edition"
// CREATED		"Sun Oct 29 11:23:20 2017"

module DIVSixteen(
	D,
	Q,
	R
);


input wire	[15:0] D;
output wire	[13:0] Q;
output wire	[2:0] R;

wire	[13:0] Q_ALTERA_SYNTHESIZED;
wire	[2:0] R_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_82;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_83;
wire	SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_85;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_73;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_77;

assign	SYNTHESIZED_WIRE_6 = 0;
assign	SYNTHESIZED_WIRE_8 = 0;
assign	SYNTHESIZED_WIRE_40 = 0;
assign	SYNTHESIZED_WIRE_42 = 0;
assign	SYNTHESIZED_WIRE_43 = 0;
assign	SYNTHESIZED_WIRE_45 = 0;
assign	SYNTHESIZED_WIRE_47 = 0;
assign	SYNTHESIZED_WIRE_49 = 0;
assign	SYNTHESIZED_WIRE_51 = 0;
assign	SYNTHESIZED_WIRE_53 = 0;
assign	SYNTHESIZED_WIRE_64 = 0;
assign	SYNTHESIZED_WIRE_66 = 0;




DIVFIVEnew	b2v_inst(
	.C(D[9]),
	.A(D[11]),
	.B(D[10]),
	.D(D[8]),
	.Q0(SYNTHESIZED_WIRE_62),
	.Q1(SYNTHESIZED_WIRE_59));


DIVFIVEnew	b2v_inst1(
	.C(D[13]),
	.A(D[15]),
	.B(D[14]),
	.D(D[12]),
	.Q0(SYNTHESIZED_WIRE_68),
	.Q1(SYNTHESIZED_WIRE_67));




DIVFIVEnew	b2v_inst12(
	.C(D[1]),
	.A(D[3]),
	.B(D[2]),
	.D(D[0]),
	.Q0(SYNTHESIZED_WIRE_4),
	.Q1(SYNTHESIZED_WIRE_1));


MODD	b2v_inst13(
	.D(D[4]),
	.A(D[7]),
	.C(D[5]),
	.B(D[6]),
	.R0(SYNTHESIZED_WIRE_78),
	.R1(SYNTHESIZED_WIRE_79),
	.R2(SYNTHESIZED_WIRE_80));


MODD	b2v_inst14(
	.D(D[0]),
	.A(D[3]),
	.C(D[1]),
	.B(D[2]),
	.R0(SYNTHESIZED_WIRE_11),
	.R1(SYNTHESIZED_WIRE_13),
	.R2(SYNTHESIZED_WIRE_15));


RCASIX	b2v_inst15(
	.A(SYNTHESIZED_WIRE_0),
	.B(SYNTHESIZED_WIRE_1),
	.Cin(SYNTHESIZED_WIRE_2),
	.C(SYNTHESIZED_WIRE_3),
	.D(SYNTHESIZED_WIRE_4),
	.E(SYNTHESIZED_WIRE_5),
	.F(SYNTHESIZED_WIRE_6),
	.G(SYNTHESIZED_WIRE_7),
	.H(SYNTHESIZED_WIRE_8),
	.I(SYNTHESIZED_WIRE_9),
	.J(SYNTHESIZED_WIRE_10),
	.O5(SYNTHESIZED_WIRE_27),
	.O4(SYNTHESIZED_WIRE_30),
	.O3(SYNTHESIZED_WIRE_32),
	.O2(SYNTHESIZED_WIRE_34),
	.O1(SYNTHESIZED_WIRE_36),
	.O0(SYNTHESIZED_WIRE_38));


CIN	b2v_inst16(
	
	.Cin(SYNTHESIZED_WIRE_2));


MODDTWO	b2v_inst17(
	
	.E0(SYNTHESIZED_WIRE_20),
	.E1(SYNTHESIZED_WIRE_22),
	.E2(SYNTHESIZED_WIRE_24));


RCATHREE	b2v_inst18(
	.A1(SYNTHESIZED_WIRE_11),
	.A2(SYNTHESIZED_WIRE_78),
	.B1(SYNTHESIZED_WIRE_13),
	.B2(SYNTHESIZED_WIRE_79),
	.C1(SYNTHESIZED_WIRE_15),
	.C2(SYNTHESIZED_WIRE_80)
	);


REMA	b2v_inst19(
	.r0(SYNTHESIZED_WIRE_78),
	.r1(SYNTHESIZED_WIRE_79),
	.r2(SYNTHESIZED_WIRE_80),
	.m3(SYNTHESIZED_WIRE_0),
	.m2(SYNTHESIZED_WIRE_3),
	.m1(SYNTHESIZED_WIRE_5),
	.m0(SYNTHESIZED_WIRE_7));


DIVFIVEnew	b2v_inst2(
	.C(D[5]),
	.A(D[7]),
	.B(D[6]),
	.D(D[4]),
	.Q0(SYNTHESIZED_WIRE_10),
	.Q1(SYNTHESIZED_WIRE_9));




RCATHREE	b2v_inst22(
	.A1(SYNTHESIZED_WIRE_20),
	.A2(SYNTHESIZED_WIRE_81),
	.B1(SYNTHESIZED_WIRE_22),
	.B2(SYNTHESIZED_WIRE_82),
	.C1(SYNTHESIZED_WIRE_24),
	.C2(SYNTHESIZED_WIRE_83)
	);


RCAFOURTEEN	b2v_inst23(
	.A(SYNTHESIZED_WIRE_84),
	.Q13(SYNTHESIZED_WIRE_27),
	.Cin(SYNTHESIZED_WIRE_28),
	.B(SYNTHESIZED_WIRE_85),
	.Q12(SYNTHESIZED_WIRE_30),
	.C(SYNTHESIZED_WIRE_86),
	.Q11(SYNTHESIZED_WIRE_32),
	.D(SYNTHESIZED_WIRE_87),
	.Q10(SYNTHESIZED_WIRE_34),
	.E(SYNTHESIZED_WIRE_84),
	.Q9(SYNTHESIZED_WIRE_36),
	.F(SYNTHESIZED_WIRE_85),
	.Q8(SYNTHESIZED_WIRE_38),
	.G(SYNTHESIZED_WIRE_86),
	.Q7(SYNTHESIZED_WIRE_40),
	.H(SYNTHESIZED_WIRE_87),
	.Q6(SYNTHESIZED_WIRE_42),
	.I(SYNTHESIZED_WIRE_43),
	.Q5(SYNTHESIZED_WIRE_44),
	.J(SYNTHESIZED_WIRE_45),
	.Q4(SYNTHESIZED_WIRE_46),
	.K(SYNTHESIZED_WIRE_47),
	.Q3(SYNTHESIZED_WIRE_48),
	.L(SYNTHESIZED_WIRE_49),
	.Q2(SYNTHESIZED_WIRE_50),
	.M(SYNTHESIZED_WIRE_51),
	.Q1(SYNTHESIZED_WIRE_52),
	.N(SYNTHESIZED_WIRE_53),
	.Q0(SYNTHESIZED_WIRE_54),
	.O13(Q_ALTERA_SYNTHESIZED[0]),
	.O12(Q_ALTERA_SYNTHESIZED[1]),
	.O11(Q_ALTERA_SYNTHESIZED[2]),
	.O10(Q_ALTERA_SYNTHESIZED[3]),
	.O9(Q_ALTERA_SYNTHESIZED[4]),
	.O8(Q_ALTERA_SYNTHESIZED[5]),
	.O7(Q_ALTERA_SYNTHESIZED[6]),
	.O6(Q_ALTERA_SYNTHESIZED[7]),
	.O5(Q_ALTERA_SYNTHESIZED[8]),
	.O4(Q_ALTERA_SYNTHESIZED[9]),
	.O3(Q_ALTERA_SYNTHESIZED[10]),
	.O2(Q_ALTERA_SYNTHESIZED[11]),
	.O1(Q_ALTERA_SYNTHESIZED[12]),
	.O0(Q_ALTERA_SYNTHESIZED[13]));


CIN	b2v_inst24(
	
	.Cin(SYNTHESIZED_WIRE_28));


MODDTWO	b2v_inst25(
	
	.E0(SYNTHESIZED_WIRE_81),
	.E1(SYNTHESIZED_WIRE_82),
	.E2(SYNTHESIZED_WIRE_83));


REMA	b2v_inst26(
	.r0(SYNTHESIZED_WIRE_81),
	.r1(SYNTHESIZED_WIRE_82),
	.r2(SYNTHESIZED_WIRE_83),
	.m3(SYNTHESIZED_WIRE_84),
	.m2(SYNTHESIZED_WIRE_85),
	.m1(SYNTHESIZED_WIRE_86),
	.m0(SYNTHESIZED_WIRE_87));





RCASIX	b2v_inst3(
	.A(SYNTHESIZED_WIRE_58),
	.B(SYNTHESIZED_WIRE_59),
	.Cin(SYNTHESIZED_WIRE_60),
	.C(SYNTHESIZED_WIRE_61),
	.D(SYNTHESIZED_WIRE_62),
	.E(SYNTHESIZED_WIRE_63),
	.F(SYNTHESIZED_WIRE_64),
	.G(SYNTHESIZED_WIRE_65),
	.H(SYNTHESIZED_WIRE_66),
	.I(SYNTHESIZED_WIRE_67),
	.J(SYNTHESIZED_WIRE_68),
	.O5(SYNTHESIZED_WIRE_44),
	.O4(SYNTHESIZED_WIRE_46),
	.O3(SYNTHESIZED_WIRE_48),
	.O2(SYNTHESIZED_WIRE_50),
	.O1(SYNTHESIZED_WIRE_52),
	.O0(SYNTHESIZED_WIRE_54));







MODDTWO	b2v_inst35(
	
	.E0(R_ALTERA_SYNTHESIZED[0]),
	.E1(R_ALTERA_SYNTHESIZED[1]),
	.E2(R_ALTERA_SYNTHESIZED[2]));


MODD	b2v_inst4(
	.D(D[12]),
	.A(D[15]),
	.C(D[13]),
	.B(D[14]),
	.R0(SYNTHESIZED_WIRE_88),
	.R1(SYNTHESIZED_WIRE_89),
	.R2(SYNTHESIZED_WIRE_90));


MODD	b2v_inst5(
	.D(D[8]),
	.A(D[11]),
	.C(D[9]),
	.B(D[10]),
	.R0(SYNTHESIZED_WIRE_73),
	.R1(SYNTHESIZED_WIRE_75),
	.R2(SYNTHESIZED_WIRE_77));


CIN	b2v_inst6(
	
	.Cin(SYNTHESIZED_WIRE_60));


REMA	b2v_inst8(
	.r0(SYNTHESIZED_WIRE_88),
	.r1(SYNTHESIZED_WIRE_89),
	.r2(SYNTHESIZED_WIRE_90),
	.m3(SYNTHESIZED_WIRE_58),
	.m2(SYNTHESIZED_WIRE_61),
	.m1(SYNTHESIZED_WIRE_63),
	.m0(SYNTHESIZED_WIRE_65));


RCATHREE	b2v_inst9(
	.A1(SYNTHESIZED_WIRE_88),
	.A2(SYNTHESIZED_WIRE_73),
	.B1(SYNTHESIZED_WIRE_89),
	.B2(SYNTHESIZED_WIRE_75),
	.C1(SYNTHESIZED_WIRE_90),
	.C2(SYNTHESIZED_WIRE_77)
	);

assign	Q = Q_ALTERA_SYNTHESIZED;
assign	R = R_ALTERA_SYNTHESIZED;

endmodule
