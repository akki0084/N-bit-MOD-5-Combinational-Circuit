-- Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus II License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 15.0.0 Build 145 04/22/2015 SJ Web Edition"
-- CREATED		"Sat Oct 28 21:27:53 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY DIV IS 
	PORT
	(
		D :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		Q :  OUT  STD_LOGIC_VECTOR(13 DOWNTO 0);
		R :  OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	);
END DIV;

ARCHITECTURE bdf_type OF DIV IS 

COMPONENT divfivenew
	PORT(C : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 Q0 : OUT STD_LOGIC;
		 Q1 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT modd
	PORT(D : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 R0 : OUT STD_LOGIC;
		 R1 : OUT STD_LOGIC;
		 R2 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT rcasix
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 E : IN STD_LOGIC;
		 F : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 H : IN STD_LOGIC;
		 I : IN STD_LOGIC;
		 J : IN STD_LOGIC;
		 O5 : OUT STD_LOGIC;
		 O4 : OUT STD_LOGIC;
		 O3 : OUT STD_LOGIC;
		 O2 : OUT STD_LOGIC;
		 O1 : OUT STD_LOGIC;
		 O0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT cin
	PORT(I : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 Cin : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT rcathree
	PORT(A1 : IN STD_LOGIC;
		 A2 : IN STD_LOGIC;
		 B1 : IN STD_LOGIC;
		 B2 : IN STD_LOGIC;
		 C1 : IN STD_LOGIC;
		 C2 : IN STD_LOGIC;
		 S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT rema
	PORT(r0 : IN STD_LOGIC;
		 r1 : IN STD_LOGIC;
		 r2 : IN STD_LOGIC;
		 m3 : OUT STD_LOGIC;
		 m2 : OUT STD_LOGIC;
		 m1 : OUT STD_LOGIC;
		 m0 : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT rcafourteen
	PORT(A : IN STD_LOGIC;
		 Q13 : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Q12 : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 Q11 : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 Q10 : IN STD_LOGIC;
		 E : IN STD_LOGIC;
		 Q9 : IN STD_LOGIC;
		 F : IN STD_LOGIC;
		 Q8 : IN STD_LOGIC;
		 G : IN STD_LOGIC;
		 Q7 : IN STD_LOGIC;
		 H : IN STD_LOGIC;
		 Q6 : IN STD_LOGIC;
		 I : IN STD_LOGIC;
		 Q5 : IN STD_LOGIC;
		 J : IN STD_LOGIC;
		 Q4 : IN STD_LOGIC;
		 K : IN STD_LOGIC;
		 Q3 : IN STD_LOGIC;
		 L : IN STD_LOGIC;
		 Q2 : IN STD_LOGIC;
		 M : IN STD_LOGIC;
		 Q1 : IN STD_LOGIC;
		 N : IN STD_LOGIC;
		 Q0 : IN STD_LOGIC;
		 O13 : OUT STD_LOGIC;
		 O12 : OUT STD_LOGIC;
		 O11 : OUT STD_LOGIC;
		 O10 : OUT STD_LOGIC;
		 O9 : OUT STD_LOGIC;
		 O8 : OUT STD_LOGIC;
		 O7 : OUT STD_LOGIC;
		 O6 : OUT STD_LOGIC;
		 O5 : OUT STD_LOGIC;
		 O4 : OUT STD_LOGIC;
		 O3 : OUT STD_LOGIC;
		 O2 : OUT STD_LOGIC;
		 O1 : OUT STD_LOGIC;
		 O0 : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	Q_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL	R_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_55 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_105 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_6 <= '0';
SYNTHESIZED_WIRE_8 <= '0';
SYNTHESIZED_WIRE_44 <= '0';
SYNTHESIZED_WIRE_46 <= '0';
SYNTHESIZED_WIRE_47 <= '0';
SYNTHESIZED_WIRE_49 <= '0';
SYNTHESIZED_WIRE_51 <= '0';
SYNTHESIZED_WIRE_53 <= '0';
SYNTHESIZED_WIRE_55 <= '0';
SYNTHESIZED_WIRE_57 <= '0';
SYNTHESIZED_WIRE_72 <= '0';
SYNTHESIZED_WIRE_74 <= '0';



b2v_inst : divfivenew
PORT MAP(C => D(9),
		 A => D(11),
		 B => D(10),
		 D => D(8),
		 Q0 => SYNTHESIZED_WIRE_70,
		 Q1 => SYNTHESIZED_WIRE_67);


b2v_inst1 : divfivenew
PORT MAP(C => D(13),
		 A => D(15),
		 B => D(14),
		 D => D(12),
		 Q0 => SYNTHESIZED_WIRE_76,
		 Q1 => SYNTHESIZED_WIRE_75);




b2v_inst12 : divfivenew
PORT MAP(C => D(1),
		 A => D(3),
		 B => D(2),
		 D => D(0),
		 Q0 => SYNTHESIZED_WIRE_4,
		 Q1 => SYNTHESIZED_WIRE_1);


b2v_inst13 : modd
PORT MAP(D => D(4),
		 A => D(7),
		 C => D(5),
		 B => D(6),
		 R0 => SYNTHESIZED_WIRE_91,
		 R1 => SYNTHESIZED_WIRE_92,
		 R2 => SYNTHESIZED_WIRE_93);


b2v_inst14 : modd
PORT MAP(D => D(0),
		 A => D(3),
		 C => D(1),
		 B => D(2),
		 R0 => SYNTHESIZED_WIRE_15,
		 R1 => SYNTHESIZED_WIRE_17,
		 R2 => SYNTHESIZED_WIRE_19);


b2v_inst15 : rcasix
PORT MAP(A => SYNTHESIZED_WIRE_0,
		 B => SYNTHESIZED_WIRE_1,
		 Cin => SYNTHESIZED_WIRE_2,
		 C => SYNTHESIZED_WIRE_3,
		 D => SYNTHESIZED_WIRE_4,
		 E => SYNTHESIZED_WIRE_5,
		 F => SYNTHESIZED_WIRE_6,
		 G => SYNTHESIZED_WIRE_7,
		 H => SYNTHESIZED_WIRE_8,
		 I => SYNTHESIZED_WIRE_9,
		 J => SYNTHESIZED_WIRE_10,
		 O5 => SYNTHESIZED_WIRE_31,
		 O4 => SYNTHESIZED_WIRE_34,
		 O3 => SYNTHESIZED_WIRE_36,
		 O2 => SYNTHESIZED_WIRE_38,
		 O1 => SYNTHESIZED_WIRE_40,
		 O0 => SYNTHESIZED_WIRE_42);


b2v_inst16 : cin
PORT MAP(		 Cin => SYNTHESIZED_WIRE_2);


b2v_inst17 : modd
PORT MAP(D => SYNTHESIZED_WIRE_90,
		 A => SYNTHESIZED_WIRE_90,
		 C => SYNTHESIZED_WIRE_90,
		 B => SYNTHESIZED_WIRE_90,
		 R0 => SYNTHESIZED_WIRE_24,
		 R1 => SYNTHESIZED_WIRE_26,
		 R2 => SYNTHESIZED_WIRE_28);


b2v_inst18 : rcathree
PORT MAP(A1 => SYNTHESIZED_WIRE_15,
		 A2 => SYNTHESIZED_WIRE_91,
		 B1 => SYNTHESIZED_WIRE_17,
		 B2 => SYNTHESIZED_WIRE_92,
		 C1 => SYNTHESIZED_WIRE_19,
		 C2 => SYNTHESIZED_WIRE_93,
		 S => SYNTHESIZED_WIRE_90);


b2v_inst19 : rema
PORT MAP(r0 => SYNTHESIZED_WIRE_91,
		 r1 => SYNTHESIZED_WIRE_92,
		 r2 => SYNTHESIZED_WIRE_93,
		 m3 => SYNTHESIZED_WIRE_0,
		 m2 => SYNTHESIZED_WIRE_3,
		 m1 => SYNTHESIZED_WIRE_5,
		 m0 => SYNTHESIZED_WIRE_7);


b2v_inst2 : divfivenew
PORT MAP(C => D(5),
		 A => D(7),
		 B => D(6),
		 D => D(4),
		 Q0 => SYNTHESIZED_WIRE_10,
		 Q1 => SYNTHESIZED_WIRE_9);




b2v_inst22 : rcathree
PORT MAP(A1 => SYNTHESIZED_WIRE_24,
		 A2 => SYNTHESIZED_WIRE_94,
		 B1 => SYNTHESIZED_WIRE_26,
		 B2 => SYNTHESIZED_WIRE_95,
		 C1 => SYNTHESIZED_WIRE_28,
		 C2 => SYNTHESIZED_WIRE_96,
		 S => SYNTHESIZED_WIRE_101);


b2v_inst23 : rcafourteen
PORT MAP(A => SYNTHESIZED_WIRE_97,
		 Q13 => SYNTHESIZED_WIRE_31,
		 Cin => SYNTHESIZED_WIRE_32,
		 B => SYNTHESIZED_WIRE_98,
		 Q12 => SYNTHESIZED_WIRE_34,
		 C => SYNTHESIZED_WIRE_99,
		 Q11 => SYNTHESIZED_WIRE_36,
		 D => SYNTHESIZED_WIRE_100,
		 Q10 => SYNTHESIZED_WIRE_38,
		 E => SYNTHESIZED_WIRE_97,
		 Q9 => SYNTHESIZED_WIRE_40,
		 F => SYNTHESIZED_WIRE_98,
		 Q8 => SYNTHESIZED_WIRE_42,
		 G => SYNTHESIZED_WIRE_99,
		 Q7 => SYNTHESIZED_WIRE_44,
		 H => SYNTHESIZED_WIRE_100,
		 Q6 => SYNTHESIZED_WIRE_46,
		 I => SYNTHESIZED_WIRE_47,
		 Q5 => SYNTHESIZED_WIRE_48,
		 J => SYNTHESIZED_WIRE_49,
		 Q4 => SYNTHESIZED_WIRE_50,
		 K => SYNTHESIZED_WIRE_51,
		 Q3 => SYNTHESIZED_WIRE_52,
		 L => SYNTHESIZED_WIRE_53,
		 Q2 => SYNTHESIZED_WIRE_54,
		 M => SYNTHESIZED_WIRE_55,
		 Q1 => SYNTHESIZED_WIRE_56,
		 N => SYNTHESIZED_WIRE_57,
		 Q0 => SYNTHESIZED_WIRE_58,
		 O13 => Q_ALTERA_SYNTHESIZED(0),
		 O12 => Q_ALTERA_SYNTHESIZED(1),
		 O11 => Q_ALTERA_SYNTHESIZED(2),
		 O10 => Q_ALTERA_SYNTHESIZED(3),
		 O9 => Q_ALTERA_SYNTHESIZED(4),
		 O8 => Q_ALTERA_SYNTHESIZED(5),
		 O7 => Q_ALTERA_SYNTHESIZED(6),
		 O6 => Q_ALTERA_SYNTHESIZED(7),
		 O5 => Q_ALTERA_SYNTHESIZED(8),
		 O4 => Q_ALTERA_SYNTHESIZED(9),
		 O3 => Q_ALTERA_SYNTHESIZED(10),
		 O2 => Q_ALTERA_SYNTHESIZED(11),
		 O1 => Q_ALTERA_SYNTHESIZED(12),
		 O0 => Q_ALTERA_SYNTHESIZED(13));


b2v_inst24 : cin
PORT MAP(		 Cin => SYNTHESIZED_WIRE_32);


b2v_inst25 : modd
PORT MAP(D => SYNTHESIZED_WIRE_101,
		 A => SYNTHESIZED_WIRE_101,
		 C => SYNTHESIZED_WIRE_101,
		 B => SYNTHESIZED_WIRE_101,
		 R0 => R_ALTERA_SYNTHESIZED(0),
		 R1 => R_ALTERA_SYNTHESIZED(1),
		 R2 => R_ALTERA_SYNTHESIZED(2));


b2v_inst26 : rema
PORT MAP(r0 => SYNTHESIZED_WIRE_94,
		 r1 => SYNTHESIZED_WIRE_95,
		 r2 => SYNTHESIZED_WIRE_96,
		 m3 => SYNTHESIZED_WIRE_97,
		 m2 => SYNTHESIZED_WIRE_98,
		 m1 => SYNTHESIZED_WIRE_99,
		 m0 => SYNTHESIZED_WIRE_100);





b2v_inst3 : rcasix
PORT MAP(A => SYNTHESIZED_WIRE_66,
		 B => SYNTHESIZED_WIRE_67,
		 Cin => SYNTHESIZED_WIRE_68,
		 C => SYNTHESIZED_WIRE_69,
		 D => SYNTHESIZED_WIRE_70,
		 E => SYNTHESIZED_WIRE_71,
		 F => SYNTHESIZED_WIRE_72,
		 G => SYNTHESIZED_WIRE_73,
		 H => SYNTHESIZED_WIRE_74,
		 I => SYNTHESIZED_WIRE_75,
		 J => SYNTHESIZED_WIRE_76,
		 O5 => SYNTHESIZED_WIRE_48,
		 O4 => SYNTHESIZED_WIRE_50,
		 O3 => SYNTHESIZED_WIRE_52,
		 O2 => SYNTHESIZED_WIRE_54,
		 O1 => SYNTHESIZED_WIRE_56,
		 O0 => SYNTHESIZED_WIRE_58);







b2v_inst4 : modd
PORT MAP(D => D(12),
		 A => D(15),
		 C => D(13),
		 B => D(14),
		 R0 => SYNTHESIZED_WIRE_103,
		 R1 => SYNTHESIZED_WIRE_104,
		 R2 => SYNTHESIZED_WIRE_105);


b2v_inst5 : modd
PORT MAP(D => D(8),
		 A => D(11),
		 C => D(9),
		 B => D(10),
		 R0 => SYNTHESIZED_WIRE_85,
		 R1 => SYNTHESIZED_WIRE_87,
		 R2 => SYNTHESIZED_WIRE_89);


b2v_inst6 : cin
PORT MAP(		 Cin => SYNTHESIZED_WIRE_68);


b2v_inst7 : modd
PORT MAP(D => SYNTHESIZED_WIRE_102,
		 A => SYNTHESIZED_WIRE_102,
		 C => SYNTHESIZED_WIRE_102,
		 B => SYNTHESIZED_WIRE_102,
		 R0 => SYNTHESIZED_WIRE_94,
		 R1 => SYNTHESIZED_WIRE_95,
		 R2 => SYNTHESIZED_WIRE_96);


b2v_inst8 : rema
PORT MAP(r0 => SYNTHESIZED_WIRE_103,
		 r1 => SYNTHESIZED_WIRE_104,
		 r2 => SYNTHESIZED_WIRE_105,
		 m3 => SYNTHESIZED_WIRE_66,
		 m2 => SYNTHESIZED_WIRE_69,
		 m1 => SYNTHESIZED_WIRE_71,
		 m0 => SYNTHESIZED_WIRE_73);


b2v_inst9 : rcathree
PORT MAP(A1 => SYNTHESIZED_WIRE_103,
		 A2 => SYNTHESIZED_WIRE_85,
		 B1 => SYNTHESIZED_WIRE_104,
		 B2 => SYNTHESIZED_WIRE_87,
		 C1 => SYNTHESIZED_WIRE_105,
		 C2 => SYNTHESIZED_WIRE_89,
		 S => SYNTHESIZED_WIRE_102);

Q <= Q_ALTERA_SYNTHESIZED;
R <= R_ALTERA_SYNTHESIZED;

END bdf_type;